BLUE
100 100 100 100 100 g c 0 1 39 1
10 10 10 10 10 g c 4 1 32 1 
10 10 10 10 10 g c 8 1 27 1 
10 10 10 10 10 g c 15 1 20 1 
4 3 0 8 4 11 3 9 1 8 1 3 5 1 4 9 3 5 0 10 3 4 2 2 1 6 1 6 2 11 0 12 0 4 2 5 2 10 
Geese is at: 12
