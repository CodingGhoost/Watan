RED
1 1 0 2 0 g 38 c 25 1 37 1 
3 1 0 0 5 g 23 c 15 1 28 1 
2 1 0 0 2 g 14 10 c 14 1 40 2 
1 0 1 0 0 g c 6 1 53 1 
1 6 4 5 1 10 2 2 0 3 1 3 3 6 4 8 3 10 0 11 0 9 0 12 4 4 2 9 5 1 1 5 2 11 3 8 2 4 
Geese is at: -1
